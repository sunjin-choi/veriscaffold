

module hello_world;
  initial begin
    $display("Hello, World from SystemVerilog!");
    $finish;
  end
endmodule
