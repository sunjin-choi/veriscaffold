// General parameterizable N x M xbar
// TODO: duplicate of selector_if?

interface xbar_if #(
    parameter type DATA_TYPE,
    parameter int  ENTRIES_X,
    parameter int  ENTRIES_Y
);

endinterface
