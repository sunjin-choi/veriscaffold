

module hello;
  initial begin
    $display("Hello, World from SystemVerilog!");
    $finish;
  end
endmodule
